module BIT_AND (Reg1, Reg2, Out);

input [15:0] Reg1, Reg2;
output [15:0] Out;

assign Out = Reg1 & Reg2;

endmodule