module NOP ();
endmodule