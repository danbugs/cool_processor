
module MOV_n (in, out);

output [15:0] out;
input [6:0] in;

assign out = in;

endmodule