module MOV (Reg1, Reg2);

input [15:0] Reg1, Reg2;

assign Reg1 = Reg2;

endmodule
