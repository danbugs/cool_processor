module ADR (Reg1, n);

input [15:0] Reg1;
input [6:0] n;

assign Reg1 = n;

endmodule
